library ieee;
use ieee.std_logic_1164.all;
package Flipflops is 
	component dff_set is port(
									  D		:in std_logic;
									  clk    :in std_logic;
									  set    :in std_logic;
									  Q      :out std_logic
									  );
	end component dff_set;
	
	component dff_reset	is port(
									  D		:in std_logic;
									  clk    :in std_logic;
									  reset  :in std_logic;
									  Q      :out std_logic
									  );
	end component dff_reset;
  
end package Flipflops;

library ieee;
use ieee.std_logic_1164.all;
	entity dff_set	is port(
								D		 :in std_logic;
								clk    :in std_logic;
								set    :in std_logic;
								Q      :out std_logic
								);
	end entity dff_set;

architecture struct of dff_set is  
begin
dff_set_proc: process (clk,set)
begin
	if(set='1')then
	Q <= '1';
	elsif (clk'event and (clk='1')) then
	Q <=D;
	end if;
	
end process dff_set_proc;
end struct;





library ieee;
use ieee.std_logic_1164.all;
entity dff_reset	is port(
									  D		:in std_logic;
									  clk	   :in std_logic;
									  reset  :in std_logic;
									  Q      :out std_logic
									  );
end entity dff_reset;

architecture struct of dff_reset is  
begin
dff_reset_proc: process (clk,reset)
begin
	if(reset='1')then
	Q <= '0';
	elsif (clk'event and (clk='1')) then
	Q <=D;
	end if;
	
end process dff_reset_proc;
end struct;